`include "transaction.sv" 
`include "generator.sv"
`include "interface.sv"
`include "driver.sv"
`include "environment.sv"
`include "program.sv"
`include "parking_system.sv"
`include "tb_top.sv"
`include "cover_properties.sv"
\\`include "cover_properties_class.sv"
\\`include "assertions.sv"
\\`include "assertions_class.sv"