interface intf(input logic clk,reset_n);
logic sensor_entrance;
logic sensor_exit;
logic [1:0] password_1;
logic [1:0] password_2;
logic GREEN_LED;
logic RED_LED;
logic [6:0] HEX_1;
logic [6:0] HEX_2;

endinterface
